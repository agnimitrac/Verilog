module state1 (
    input 
);

endmodule