module moduleName #(
    parameters
) (
    ports
);
    
endmodule

module moduleName (
    ports
);
    
endmodule