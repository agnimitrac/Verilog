module tb;
    test dut();
endmodule